// qsys.v

// Generated using ACDS version 13.1 162 at 2023.12.18.02:35:13

`timescale 1 ps / 1 ps
module qsys (
		input  wire        clk_50m_clk,      //   clk_50m.clk
		input  wire        reset_reset_n,    //     reset.reset_n
		input  wire        areset_export,    //    areset.export
		output wire        locked_export,    //    locked.export
		output wire        phasedone_export, // phasedone.export
		output wire [11:0] sdram_addr,       //     sdram.addr
		output wire [1:0]  sdram_ba,         //          .ba
		output wire        sdram_cas_n,      //          .cas_n
		output wire        sdram_cke,        //          .cke
		output wire        sdram_cs_n,       //          .cs_n
		inout  wire [15:0] sdram_dq,         //          .dq
		output wire [1:0]  sdram_dqm,        //          .dqm
		output wire        sdram_ras_n,      //          .ras_n
		output wire        sdram_we_n,       //          .we_n
		output wire        sdram_clk_clk     // sdram_clk.clk
	);

	wire         pll_c0_clk;                                                // pll:c0 -> [apb:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, mm_interconnect_0:pll_c0_clk, mm_interconnect_1:pll_c0_clk, nios2cpu:clk, rst_controller_001:clk, sdram:clk]
	wire         pll_c2_clk;                                                // pll:c2 -> [floor_timer:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, jtag_uart:clk, mm_interconnect_1:pll_c2_clk, rst_controller_002:clk, seg7_timer:clk, sys_timer:clk]
	wire         nios2cpu_instruction_master_waitrequest;                   // mm_interconnect_0:nios2cpu_instruction_master_waitrequest -> nios2cpu:i_waitrequest
	wire  [25:0] nios2cpu_instruction_master_address;                       // nios2cpu:i_address -> mm_interconnect_0:nios2cpu_instruction_master_address
	wire         nios2cpu_instruction_master_read;                          // nios2cpu:i_read -> mm_interconnect_0:nios2cpu_instruction_master_read
	wire  [31:0] nios2cpu_instruction_master_readdata;                      // mm_interconnect_0:nios2cpu_instruction_master_readdata -> nios2cpu:i_readdata
	wire         mm_interconnect_0_apb_s0_waitrequest;                      // apb:s0_waitrequest -> mm_interconnect_0:apb_s0_waitrequest
	wire   [0:0] mm_interconnect_0_apb_s0_burstcount;                       // mm_interconnect_0:apb_s0_burstcount -> apb:s0_burstcount
	wire  [31:0] mm_interconnect_0_apb_s0_writedata;                        // mm_interconnect_0:apb_s0_writedata -> apb:s0_writedata
	wire   [9:0] mm_interconnect_0_apb_s0_address;                          // mm_interconnect_0:apb_s0_address -> apb:s0_address
	wire         mm_interconnect_0_apb_s0_write;                            // mm_interconnect_0:apb_s0_write -> apb:s0_write
	wire         mm_interconnect_0_apb_s0_read;                             // mm_interconnect_0:apb_s0_read -> apb:s0_read
	wire  [31:0] mm_interconnect_0_apb_s0_readdata;                         // apb:s0_readdata -> mm_interconnect_0:apb_s0_readdata
	wire         mm_interconnect_0_apb_s0_debugaccess;                      // mm_interconnect_0:apb_s0_debugaccess -> apb:s0_debugaccess
	wire         mm_interconnect_0_apb_s0_readdatavalid;                    // apb:s0_readdatavalid -> mm_interconnect_0:apb_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_apb_s0_byteenable;                       // mm_interconnect_0:apb_s0_byteenable -> apb:s0_byteenable
	wire         nios2cpu_data_master_waitrequest;                          // mm_interconnect_0:nios2cpu_data_master_waitrequest -> nios2cpu:d_waitrequest
	wire  [31:0] nios2cpu_data_master_writedata;                            // nios2cpu:d_writedata -> mm_interconnect_0:nios2cpu_data_master_writedata
	wire  [25:0] nios2cpu_data_master_address;                              // nios2cpu:d_address -> mm_interconnect_0:nios2cpu_data_master_address
	wire         nios2cpu_data_master_write;                                // nios2cpu:d_write -> mm_interconnect_0:nios2cpu_data_master_write
	wire         nios2cpu_data_master_read;                                 // nios2cpu:d_read -> mm_interconnect_0:nios2cpu_data_master_read
	wire  [31:0] nios2cpu_data_master_readdata;                             // mm_interconnect_0:nios2cpu_data_master_readdata -> nios2cpu:d_readdata
	wire         nios2cpu_data_master_debugaccess;                          // nios2cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2cpu_data_master_debugaccess
	wire   [3:0] nios2cpu_data_master_byteenable;                           // nios2cpu:d_byteenable -> mm_interconnect_0:nios2cpu_data_master_byteenable
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                 // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                   // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_write;                     // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_0_pll_pll_slave_read;                      // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                  // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_nios2cpu_jtag_debug_module_waitrequest;  // nios2cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2cpu_jtag_debug_module_writedata;    // mm_interconnect_0:nios2cpu_jtag_debug_module_writedata -> nios2cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2cpu_jtag_debug_module_address;      // mm_interconnect_0:nios2cpu_jtag_debug_module_address -> nios2cpu:jtag_debug_module_address
	wire         mm_interconnect_0_nios2cpu_jtag_debug_module_write;        // mm_interconnect_0:nios2cpu_jtag_debug_module_write -> nios2cpu:jtag_debug_module_write
	wire         mm_interconnect_0_nios2cpu_jtag_debug_module_read;         // mm_interconnect_0:nios2cpu_jtag_debug_module_read -> nios2cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2cpu_jtag_debug_module_readdata;     // nios2cpu:jtag_debug_module_readdata -> mm_interconnect_0:nios2cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2cpu_jtag_debug_module_debugaccess;  // mm_interconnect_0:nios2cpu_jtag_debug_module_debugaccess -> nios2cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2cpu_jtag_debug_module_byteenable;   // mm_interconnect_0:nios2cpu_jtag_debug_module_byteenable -> nios2cpu:jtag_debug_module_byteenable
	wire   [0:0] apb_m0_burstcount;                                         // apb:m0_burstcount -> mm_interconnect_1:apb_m0_burstcount
	wire         apb_m0_waitrequest;                                        // mm_interconnect_1:apb_m0_waitrequest -> apb:m0_waitrequest
	wire   [9:0] apb_m0_address;                                            // apb:m0_address -> mm_interconnect_1:apb_m0_address
	wire  [31:0] apb_m0_writedata;                                          // apb:m0_writedata -> mm_interconnect_1:apb_m0_writedata
	wire         apb_m0_write;                                              // apb:m0_write -> mm_interconnect_1:apb_m0_write
	wire         apb_m0_read;                                               // apb:m0_read -> mm_interconnect_1:apb_m0_read
	wire  [31:0] apb_m0_readdata;                                           // mm_interconnect_1:apb_m0_readdata -> apb:m0_readdata
	wire         apb_m0_debugaccess;                                        // apb:m0_debugaccess -> mm_interconnect_1:apb_m0_debugaccess
	wire   [3:0] apb_m0_byteenable;                                         // apb:m0_byteenable -> mm_interconnect_1:apb_m0_byteenable
	wire         apb_m0_readdatavalid;                                      // mm_interconnect_1:apb_m0_readdatavalid -> apb:m0_readdatavalid
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_1_sys_timer_s1_writedata;                  // mm_interconnect_1:sys_timer_s1_writedata -> sys_timer:writedata
	wire   [2:0] mm_interconnect_1_sys_timer_s1_address;                    // mm_interconnect_1:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_1_sys_timer_s1_chipselect;                 // mm_interconnect_1:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire         mm_interconnect_1_sys_timer_s1_write;                      // mm_interconnect_1:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_timer_s1_readdata;                   // sys_timer:readdata -> mm_interconnect_1:sys_timer_s1_readdata
	wire  [15:0] mm_interconnect_1_seg7_timer_s1_writedata;                 // mm_interconnect_1:seg7_timer_s1_writedata -> seg7_timer:writedata
	wire   [2:0] mm_interconnect_1_seg7_timer_s1_address;                   // mm_interconnect_1:seg7_timer_s1_address -> seg7_timer:address
	wire         mm_interconnect_1_seg7_timer_s1_chipselect;                // mm_interconnect_1:seg7_timer_s1_chipselect -> seg7_timer:chipselect
	wire         mm_interconnect_1_seg7_timer_s1_write;                     // mm_interconnect_1:seg7_timer_s1_write -> seg7_timer:write_n
	wire  [15:0] mm_interconnect_1_seg7_timer_s1_readdata;                  // seg7_timer:readdata -> mm_interconnect_1:seg7_timer_s1_readdata
	wire  [15:0] mm_interconnect_1_floor_timer_s1_writedata;                // mm_interconnect_1:floor_timer_s1_writedata -> floor_timer:writedata
	wire   [2:0] mm_interconnect_1_floor_timer_s1_address;                  // mm_interconnect_1:floor_timer_s1_address -> floor_timer:address
	wire         mm_interconnect_1_floor_timer_s1_chipselect;               // mm_interconnect_1:floor_timer_s1_chipselect -> floor_timer:chipselect
	wire         mm_interconnect_1_floor_timer_s1_write;                    // mm_interconnect_1:floor_timer_s1_write -> floor_timer:write_n
	wire  [15:0] mm_interconnect_1_floor_timer_s1_readdata;                 // floor_timer:readdata -> mm_interconnect_1:floor_timer_s1_readdata
	wire  [31:0] nios2cpu_d_irq_irq;                                        // irq_mapper:sender_irq -> nios2cpu:d_irq
	wire         irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                         // sys_timer:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                  // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                         // floor_timer:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                  // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                         // seg7_timer:irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [apb:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_interconnect_0:nios2cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:apb_reset_reset_bridge_in_reset_reset, nios2cpu:reset_n, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios2cpu:reset_req, rst_translator:reset_req_in]
	wire         nios2cpu_jtag_debug_module_reset_reset;                    // nios2cpu:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [floor_timer:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart:rst_n, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, seg7_timer:reset_n, sys_timer:reset_n]

	qsys_pll pll (
		.clk       (clk_50m_clk),                               //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (sdram_clk_clk),                             //                    c1.clk
		.c2        (pll_c2_clk),                                //                    c2.clk
		.areset    (areset_export),                             //        areset_conduit.export
		.locked    (locked_export),                             //        locked_conduit.export
		.phasedone (phasedone_export)                           //     phasedone_conduit.export
	);

	qsys_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	qsys_nios2cpu nios2cpu (
		.clk                                   (pll_c0_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (nios2cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2cpu_data_master_read),                                //                          .read
		.d_readdata                            (nios2cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2cpu_data_master_write),                               //                          .write
		.d_writedata                           (nios2cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                          // custom_instruction_master.readra
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) apb (
		.clk              (pll_c0_clk),                             //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),     // reset.reset
		.s0_waitrequest   (mm_interconnect_0_apb_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_apb_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_apb_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_apb_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_apb_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_apb_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_apb_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_apb_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_apb_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_apb_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (apb_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (apb_m0_readdata),                        //      .readdata
		.m0_readdatavalid (apb_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (apb_m0_burstcount),                      //      .burstcount
		.m0_writedata     (apb_m0_writedata),                       //      .writedata
		.m0_address       (apb_m0_address),                         //      .address
		.m0_write         (apb_m0_write),                           //      .write
		.m0_read          (apb_m0_read),                            //      .read
		.m0_byteenable    (apb_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (apb_m0_debugaccess)                      //      .debugaccess
	);

	qsys_jtag_uart jtag_uart (
		.clk            (pll_c2_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                              //               irq.irq
	);

	qsys_sys_timer sys_timer (
		.clk        (pll_c2_clk),                                //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)          //   irq.irq
	);

	qsys_sys_timer floor_timer (
		.clk        (pll_c2_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_floor_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_floor_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_floor_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_floor_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_floor_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)            //   irq.irq
	);

	qsys_sys_timer seg7_timer (
		.clk        (pll_c2_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),        // reset.reset_n
		.address    (mm_interconnect_1_seg7_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_seg7_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_seg7_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_seg7_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_seg7_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_003_receiver_irq)           //   irq.irq
	);

	qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_50m_clk_clk                                       (clk_50m_clk),                                              //                                     clk_50m_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                               //                                          pll_c0.clk
		.nios2cpu_reset_n_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                       //          nios2cpu_reset_n_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2cpu_data_master_address                          (nios2cpu_data_master_address),                             //                            nios2cpu_data_master.address
		.nios2cpu_data_master_waitrequest                      (nios2cpu_data_master_waitrequest),                         //                                                .waitrequest
		.nios2cpu_data_master_byteenable                       (nios2cpu_data_master_byteenable),                          //                                                .byteenable
		.nios2cpu_data_master_read                             (nios2cpu_data_master_read),                                //                                                .read
		.nios2cpu_data_master_readdata                         (nios2cpu_data_master_readdata),                            //                                                .readdata
		.nios2cpu_data_master_write                            (nios2cpu_data_master_write),                               //                                                .write
		.nios2cpu_data_master_writedata                        (nios2cpu_data_master_writedata),                           //                                                .writedata
		.nios2cpu_data_master_debugaccess                      (nios2cpu_data_master_debugaccess),                         //                                                .debugaccess
		.nios2cpu_instruction_master_address                   (nios2cpu_instruction_master_address),                      //                     nios2cpu_instruction_master.address
		.nios2cpu_instruction_master_waitrequest               (nios2cpu_instruction_master_waitrequest),                  //                                                .waitrequest
		.nios2cpu_instruction_master_read                      (nios2cpu_instruction_master_read),                         //                                                .read
		.nios2cpu_instruction_master_readdata                  (nios2cpu_instruction_master_readdata),                     //                                                .readdata
		.apb_s0_address                                        (mm_interconnect_0_apb_s0_address),                         //                                          apb_s0.address
		.apb_s0_write                                          (mm_interconnect_0_apb_s0_write),                           //                                                .write
		.apb_s0_read                                           (mm_interconnect_0_apb_s0_read),                            //                                                .read
		.apb_s0_readdata                                       (mm_interconnect_0_apb_s0_readdata),                        //                                                .readdata
		.apb_s0_writedata                                      (mm_interconnect_0_apb_s0_writedata),                       //                                                .writedata
		.apb_s0_burstcount                                     (mm_interconnect_0_apb_s0_burstcount),                      //                                                .burstcount
		.apb_s0_byteenable                                     (mm_interconnect_0_apb_s0_byteenable),                      //                                                .byteenable
		.apb_s0_readdatavalid                                  (mm_interconnect_0_apb_s0_readdatavalid),                   //                                                .readdatavalid
		.apb_s0_waitrequest                                    (mm_interconnect_0_apb_s0_waitrequest),                     //                                                .waitrequest
		.apb_s0_debugaccess                                    (mm_interconnect_0_apb_s0_debugaccess),                     //                                                .debugaccess
		.nios2cpu_jtag_debug_module_address                    (mm_interconnect_0_nios2cpu_jtag_debug_module_address),     //                      nios2cpu_jtag_debug_module.address
		.nios2cpu_jtag_debug_module_write                      (mm_interconnect_0_nios2cpu_jtag_debug_module_write),       //                                                .write
		.nios2cpu_jtag_debug_module_read                       (mm_interconnect_0_nios2cpu_jtag_debug_module_read),        //                                                .read
		.nios2cpu_jtag_debug_module_readdata                   (mm_interconnect_0_nios2cpu_jtag_debug_module_readdata),    //                                                .readdata
		.nios2cpu_jtag_debug_module_writedata                  (mm_interconnect_0_nios2cpu_jtag_debug_module_writedata),   //                                                .writedata
		.nios2cpu_jtag_debug_module_byteenable                 (mm_interconnect_0_nios2cpu_jtag_debug_module_byteenable),  //                                                .byteenable
		.nios2cpu_jtag_debug_module_waitrequest                (mm_interconnect_0_nios2cpu_jtag_debug_module_waitrequest), //                                                .waitrequest
		.nios2cpu_jtag_debug_module_debugaccess                (mm_interconnect_0_nios2cpu_jtag_debug_module_debugaccess), //                                                .debugaccess
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                  //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                    //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                     //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                 //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                //                                                .writedata
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                       //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                         //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                          //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                      //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                     //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                    //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                 //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                   //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect)                     //                                                .chipselect
	);

	qsys_mm_interconnect_1 mm_interconnect_1 (
		.pll_c0_clk                                  (pll_c0_clk),                                                //                                pll_c0.clk
		.pll_c2_clk                                  (pll_c2_clk),                                                //                                pll_c2.clk
		.apb_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                        //       apb_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // jtag_uart_reset_reset_bridge_in_reset.reset
		.apb_m0_address                              (apb_m0_address),                                            //                                apb_m0.address
		.apb_m0_waitrequest                          (apb_m0_waitrequest),                                        //                                      .waitrequest
		.apb_m0_burstcount                           (apb_m0_burstcount),                                         //                                      .burstcount
		.apb_m0_byteenable                           (apb_m0_byteenable),                                         //                                      .byteenable
		.apb_m0_read                                 (apb_m0_read),                                               //                                      .read
		.apb_m0_readdata                             (apb_m0_readdata),                                           //                                      .readdata
		.apb_m0_readdatavalid                        (apb_m0_readdatavalid),                                      //                                      .readdatavalid
		.apb_m0_write                                (apb_m0_write),                                              //                                      .write
		.apb_m0_writedata                            (apb_m0_writedata),                                          //                                      .writedata
		.apb_m0_debugaccess                          (apb_m0_debugaccess),                                        //                                      .debugaccess
		.floor_timer_s1_address                      (mm_interconnect_1_floor_timer_s1_address),                  //                        floor_timer_s1.address
		.floor_timer_s1_write                        (mm_interconnect_1_floor_timer_s1_write),                    //                                      .write
		.floor_timer_s1_readdata                     (mm_interconnect_1_floor_timer_s1_readdata),                 //                                      .readdata
		.floor_timer_s1_writedata                    (mm_interconnect_1_floor_timer_s1_writedata),                //                                      .writedata
		.floor_timer_s1_chipselect                   (mm_interconnect_1_floor_timer_s1_chipselect),               //                                      .chipselect
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.seg7_timer_s1_address                       (mm_interconnect_1_seg7_timer_s1_address),                   //                         seg7_timer_s1.address
		.seg7_timer_s1_write                         (mm_interconnect_1_seg7_timer_s1_write),                     //                                      .write
		.seg7_timer_s1_readdata                      (mm_interconnect_1_seg7_timer_s1_readdata),                  //                                      .readdata
		.seg7_timer_s1_writedata                     (mm_interconnect_1_seg7_timer_s1_writedata),                 //                                      .writedata
		.seg7_timer_s1_chipselect                    (mm_interconnect_1_seg7_timer_s1_chipselect),                //                                      .chipselect
		.sys_timer_s1_address                        (mm_interconnect_1_sys_timer_s1_address),                    //                          sys_timer_s1.address
		.sys_timer_s1_write                          (mm_interconnect_1_sys_timer_s1_write),                      //                                      .write
		.sys_timer_s1_readdata                       (mm_interconnect_1_sys_timer_s1_readdata),                   //                                      .readdata
		.sys_timer_s1_writedata                      (mm_interconnect_1_sys_timer_s1_writedata),                  //                                      .writedata
		.sys_timer_s1_chipselect                     (mm_interconnect_1_sys_timer_s1_chipselect)                  //                                      .chipselect
	);

	qsys_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2cpu_d_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_50m_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (pll_c2_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
